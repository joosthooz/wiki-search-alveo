library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use work.snappy_tta_imem_mau.all;

package snappy_tta_imem_image is

  type std_logic_imem_matrix is array (natural range <>) of std_logic_vector(IMEMMAUWIDTH-1 downto 0);

  constant imem_array : std_logic_imem_matrix := (
"11111111011111111111111111111000111111111111111111111111111111001111111000000000000000000000000000000000011",
"01111111011111000000111010111000111111111111111111111111111111000100110100111111111111001001000000000111010",
"01111111011111111111111111111111000000000011111111111111111111111111111111111111111111001100000000000110100",
"00000001001111111111111111111000111111111111111111111111111111001000101000111111111111000000000001101111000",
"01111111011111111111111111111010000000000010001110001111111111000100010000111111111111000000000000000111010",
"01111111011111111111111111110000000000000111111111111111111111111111111111111111111111001100000000000110100",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111000000000001001111000",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111",
"01111111011111111111111111110000001000000111111111111111111111111111111111111111111111111111111111111111111",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111000000000001010111001",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111",
"00000110001001111111111111111000111111111111111111111111111111111111111111111111111111000000000000000111010",
"01111111011111111111111111110000000000010011111111111111111111111111111111111111111111111111111111111111111",
"01111111011111111111111111110000000000000111111111111111111111111111111111111111111111111111111111111111111",
"11111111011111111111111111111000111111111100001011001111111111000001111111000000000000000000000000000000000",
"01111111011111111111111111111000111111111111111111111111111111111111111111001000100100000000010000000100001",
"00010010101001111111111111111000111111111110001110001111111111000000010110111111111111000000011111111100001",
"01111111011111000000110001111000111111111110001100001000100100111111111111001000110100111111111111111111111",
"01111111011111111111111111111000111111111110000101111000111000000111100000111111111111010000000001111111001",
"01111111011110000011011000111101000000010011111111111000100000111111111111111111111111111111111111111111111",
"01111111011111111111111111111101000000000111111111111111111111111111111111111111111111111111111111111111111",
"00000110111001111111111111111000111111111111111111111111111111000000100001111111111111111111111111111111111",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111",
"01111111011111111111111111111000111111111111111111111111111111100000100100111111111111111111111111111111111",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111010000010101001111001",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111100000000000000000100",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111100000000000001000111",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111000000011110000000101",
"01111111011111111111111111110000000110011011111111111111111111111111111111111111111111000000000100111111001",
"01111111011111111111111111110000000000100011111111111111111111111111111111111111111111111111111111111111111",
"01111111011111111111111111110000000000100111111111111111111111111111111111111111111111111111111111111111111",
"00100110010000010101011000111101000000100011111111111111111111111111111111111111111111111111111111111111111",
"01111111011111111111111111111101000000100111111111111111111111111111111111111111111111111111111111111111111",
"00100110010110000011011000111000111111111111111111111111111111111111111111111111111111111111111111111111111",
"01111111011111111111111111111000111111111111111111111111111111100000100100111111111111111111111111111111111",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111100000010101001111001",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111",
"01111111011111111111111111111000111111111100001011001111111111111111111111111111111111111111111111111111111",
"01111111011111111111111111111100000000101011111111111111111111000011000001001000100100111111111111111111111",
"01111111011111111111111111111010000000110110001110001111111111000000010110111111111111111111111111111111111",
"01111111011111111111111111111000111111111111111111111000100100111111111111111111111111000000011111100100001",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111100000000110110111001",
"01111111011111111111111111111000111111111110001110001111111111000010011001111111111111111111111111111111111",
"00110110101001111111111111111111000000110011111111111111111111111111111111010001000110111111111111111111111",
"11111111011111111111111111111000111111111110001001001111111111000011111111000000000000000000000000000000000",
"01111111011111111111111111111000111111111100001011001111111111111111111111111111111111010000001000000111001",
"01111111011111000000110001111000111111111111111111111111111111111111111111001000110100111111111111111111111",
"00110010101001111111111111111111000000101011111111111111111111111111111111010000101000100000000111000100001",
"01111111011111111111111111111000111111111110001110001111111111000101010111111111111111111111111111111111111",
"00110011001000010101010000111000111111111111111111111000000101000111010001111111111111000000001001010111001",
"01111111011111111111111111111010000000101111111111111000110000000100100000111111111111111111111111111111111",
"01111111011111111111111111111101000000101011111111111111111111111111111111111111111111111111111111111111111",
"11111111011111111111111111111000111111111111111111111111111111000011111111000000000000000000000000000000000",
"00101011001001000000110001111000111111111111111111111111111111111111111111111111111111111111111111111111111",
"00010110111001111111111111111000111111111111111111111000100011111111111111111111111111111111111111111111111",
"01111111011111111111111111111000111111111111111111111111111111100000100100111111111111111111111111111111111",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111100000001101000111001",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111000000001111000111001",
"00110010111001111111111111111000111111111111111111111111111111000001100000111111111111111111111111111111111",
"01111111011111111111111111111101000000101011111111111111111111111111111111111111111111111111111111111111111",
"00110111001001111111111111111000111111111111111111111111111111000010010010001000100100000000011111111100001",
"01111111011111111111111111111000111111111110001110001000100100001000010111111111111111111111111111111111111",
"00101011001001111111111111111000111111111111111111111000010101111111111111111111111111010000001001010111001",
"00110010111001111111111111111111000000101111111111111111111111000001100000100000101000111111111111111111111",
"01111111011111111111111111111101000000101011111111111111111111111111111111101000100100100000011111111100001",
"11111111011111111111111111111000111111111111111111111111111111000000010000000000000000000000000000000000000",
"11111111011111000000110111111000111111111110001110000000101100000000011000000000000000000000000000000000000",
"00101110101001000000110111111000111111111111111111111000000101111111111111001000110100111111111111111111111",
"01111111011111111111111111111000111111111110000101011000111000111111111111111111111111111111111111111111111",
"01111111011111111111111111111111000000101111111111111111111111111111111111111111111111111111111111111111111",
"00101010111001111111111111111000111111111111111111111111111111011111100000111111111111111111111111111111111",
"00011010111001111111111111111000111111111111111111111111111111100000100011111111111111111111111111111111111",
"01111111011111111111111111111000111111111111111111111111111111100000100100111111111111111111111111111111111",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111010000001011001111001",
"00101011001001111111111111111000111111111111111111111111111111000011010001111111111111111111111111111111111",
"01111111011111111111111111111111000000110011111111111111111111111111111111111111111111111111111111111111111",
"00110001110100010101100000111000111111111111111111111111111111111111111111111111111111111111111111111111111",
"01111111011111111111111111111111000000110111111111111111111111111111111111111111111111111111111111111111111",
"00110111001001111111111111111000111111111111111111111111111111000100010000111111111111111111111111111111111",
"00101111000000010001100100111111000000110111111111111000110000000000100001111111111111111111111111111111111",
"00101111000001111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111",
"00101111000001111111111111011000111111111111111111111111111111100000100100111111111111111111111111111111111",
"00101111000001111111111111011000111111111111111111111111111111111111111111111111111111100000001010011111001",
"01111111011111111111111111011000111111111111111111111111111111111111111111111111111111111111111111111111111",
"00110111001001111111111111011000111111111111111111111111111111000100010000111111111111111111111111111111111",
"00110010111001111111111111111000111111111111111111111111111111000000100001111111111111111111111111111111111",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111",
"01111111011111111111111111111000111111111111111111111111111111100000100100111111111111111111111111111111111",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111010000000100000111001",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111",
"00100010111001111111111111111000111111111111111111111111111111111111111111010001100000111111111111111111111",
"00110010101001111111111111111000111111111111111111111111111111011111000000111111111111111111111111111111111",
"01111111011111111111111111111010000000110010001110001111111111000000010110111111111111111111111111111111111",
"01111111011111111111111111111000111111111111111111111000100100111111111111111111111111111111111111111111111",
"00101111000000010001100100111000111111111111111111111111111111111111111111111111111111010000001100000111001",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111",
"00110010101001111111111111011000111111111111111111111111111111111111111111010111000000111111111111111111111",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111000000000100000111001",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111",
"00100010111001111111111111111000111111111111111111111111111111000001100000111111111111111111111111111111111",
"00011100010101111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111",
"00010000010111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111",
"00101110101001111111111111111000111111111111111111111111111111111111111111111111111111000000011111111100001",
"10110010101001111111111111111010000000101111111111110111000000000011111111000000000000000000000000000000000",
"11111111011111000000110001111010000000110010001110001111111111000000111011000000000000000000000000000000000",
"11111111011111000001000011111000111111111100001011001000110000000011111111000000000000000000000000000000000",
"01111111011111000000110001111000111111111111111111111111111111100000100100001000110100111111111111111111111",
"00101110111000010110110111111000111111111111111111111000111000001000100000111111111111010000001101011111001",
"01111111011110010101011000111101000000101111111111111000100000111111111111111111111111111111111111111111111",
"00101110101001111111111111111101000000101011111111111111111111111111111111111111111111010000011111111100001",
"00101010111001111111111111111000111111111111111111111111111111000000100001111111111111111111111111111111111",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111",
"01111111011111111111111111111000111111111111111111111111111111100000100100111111111111111111111111111111111",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111010000000100011111001",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111",
"00100110010110000011011000111000111111111111111111111111111111111111111111111111111111111111111111111111111",
"00101010010000010011011000111000111111111111111111111111111111111111111111111111111111111111111111111111111",
"00100110010111111111111111111101000000101111111111111111111111100000101100111111111111111111111111111111111",
"01111111011111111111111111111000111111111111111111111111111111100000100100111111111111111111111111111111111",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111100000000100011111001",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111",
"00100110010110000011011000111000111111111111111111111111111111111111111111111111111111111111111111111111111",
"00101011001001111111111111111000111111111111111111111111111111000011010001111111111111111111111111111111111",
"01111111011111111111111111111111000000110111111111111000110000000000100001111111111111111111111111111111111",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111",
"01111111011111111111111111111000111111111111111111111111111111100000100100111111111111111111111111111111111",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111010000010001110111001",
"00101010111000010010001110111000111111111111111111111111111111011111100000111111111111111111111111111111111",
"01111111011111111111111111111101000000110011111111111111111111111111111111111111111111111111111111111111111",
"00110100011101111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111",
"00111010101001111111111111111000111111111111111111111111111111011111000000111111111111111111111111111111111",
"01111111011111111111111111111010000000111010001110001111111111000000010110111111111111111111111111111111111",
"01111111011111111111111111111000111111111111111111111000100100111111111111111111111111111111111111111111111",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111010000010000111111001",
"01111111011111111111111111111000111111111100001011001111111111111111111111111111111111111111111111111111111",
"00111010101001111111111111001000111111111111111111111111111111111111111111010111000000111111111111111111111",
"00110110010000010011011000111000111111111111111111111111111111111111111111111111111111111111111111111111111",
"01111111011111111111111111111101000000111011111111111111111111111111111111111111111111111111111111111111111",
"00110010010110001101011000111000111111111111111111111111111111111111111111111111111111111111111111111111111",
"01111111011111111111111111111000111111111111111111111111111111100000100100111111111111111111111111111111111",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111100000010011011111001",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111",
"00100110010000010101011000111000111111111111111111111111111111111111111111111111111111111111111111111111111",
"00101110010110000011011000111000111111111111111111111111111111111111111111111111111111111111111111111111111",
"01111111011111111111111111111000111111111111111111111111111111100000100100111111111111111111111111111111111",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111010000000101000111001",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111",
"00101100010011111111111111111000111111111111111111111111111111111111111111010000101000111111111111111111111",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111000000010101001111001",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111",
"00111011001001111111111111111000111111111111111111111111111111100000011010111111111111111111111111111111111",
"01111111011111111111111111111111000000100111111111111111111111111111111111111111111111111111111111111111111",
"00100111001001111111111111111000111111111111111111111111111111011100010000111111111111111111111111111111111",
"01111111011111111111111111111111000000100111111111111000110000000000100001111111111111111111111111111111111",
"01111111011111111111111111111000111111111100001011001111111111111111111111111111111111111111111111111111111",
"01111111011111111111111111001000111111111100001011001111111111100000100100111111111111111111111111111111111",
"01111111011111111111111111001000111111111100001011001111111111111111111111111111111111100000010011110111001",
"01111111011111111111111111001000111111111100001011001111111111111111111111111111111111111111111111111111111",
"00100111001001111111111111001000111111111111111111111111111111111111111111100100010000111111111111111111111",
"00101110010110000011011000111000111111111111111111111111111111111111111111111111111111111111111111111111111",
"01111111011111111111111111111000111111111111111111111111111111100000100100111111111111111111111111111111111",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111010000000101000111001",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111",
"00101100010011111111111111111000111111111111111111111111111111111111111111010000101000111111111111111111111",
"11111111011111111111111111111000111111111111111111111111111111001111111100000000000000000000000000000000011",
"01111111011111111111111111111000111111111111111111111111111111111111111111111111111111001001000000000111001",
"01111111011111111111111111111011000000000111111111111111111111111111111111111111111111111111111111111111111",
"00000110001001111111111111110000000000000111111111111111111111111111111111111111111111000000000000001111010");

end snappy_tta_imem_image;
