library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use work.snappy_tta_imem_mau.all;

package snappy_tta_imem_image is

  type std_logic_imem_matrix is array (natural range <>) of std_logic_vector(IMEMMAUWIDTH-1 downto 0);

  constant imem_array : std_logic_imem_matrix := (
"0111111100111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111",
"1111111100111000000010010011001111111111111111111111111111111111111000000000000000000000000000000000011",
"0111111100111110000000001001111111111111111111111111111111111111111111111111111110010010000000000111110",
"0111111100111000000100010101001111111111000011010111111111111111111111111111111110000000000001100111100",
"0111111100111111111111111111110111000000100100100100010110011111111111111111111110010100000000000110100",
"0111111100111000000000010001001111111111111111111111111111111111111111111111111110011000000000000110100",
"0111111100111000000000100001011111111111111111111111111111111111111111111111111110000000000010100111101",
"0111111100111001111000000001001111111111111111111111111111111111111111111111111111111111111111111111111",
"0111111100111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111",
"0111111100111111111111111111111111111110000100010111111111111111111111111111111111111111111111111111111",
"0000010000110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"0000010000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"0111111100111111111111111111111111111110000100011111111111111111111111111111111111111111111111111111111",
"0111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"0111111100111001000000001100011111111111111111111111111111111111111110010001110001111111111111111111111",
"0001111011000001111111101000011111111110000010110100011000011111111111111111111111111111111111111111111",
"0111111100111000111111101100010011001111000101100100010010011111111110010001110001111111111111111111111",
"0111111100111100000011101101111111111110111100100100011000011111111111111111111110100000000011100111101",
"0111111100111100000011010100000110001111111111111100010000011111111111111111111110100000000000000111011",
"0111111100111111111111111111110110001101111111111111111111111111111111111111111111111111111111111111111",
"0001101011100111111111111111111111111110000100101111111111111111111111111111111111111111111111111111111",
"0111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"0111111100111111111111111111111111111111111111111111111111110001001001111111111111111111111111111111111",
"0111111100111111111111111111111111111111111111111111111111111111111111111111111110100000000010100111101",
"0111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"0111111100111111111111111111111111111111111111111111111111111111111111111111111110100000000000000111010",
"0111111100111111111111111111111111111111111111111111111111111111111111111111111110000000001001110111101",
"0111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"0000010000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"0010001100000111111111111111110011010100111010001111111111111111111111111111111111111111111111111111111",
"0010101100000000000010010000001111111110101010111100010110011111111111111111111111111111111111111111111",
"0010011100000111111111111111110110010001111111111100001010111111111111111111111111111111111111111111111",
"0001111001100100000100010100000111010011111111111111111111111111111111111111111111111111111111111111111",
"0010001001001100000100110110000110001111111111111111111111111111111111111111111111111111111111111111111",
"0001111001111100000011010100001111111111111111111111111111111111111111111111111111111111111111111111111",
"0111111100111111111111111111111111111111111111111111111111110001001001111111111111111111111111111111111",
"0111111100111111111111111111111111111111111111111111111111111111111111111111111111000000000010100111101",
"0111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"0111111100111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111010",
"0111111100111111111111111111111111111110000100011111111111111111111111111111111111111111111111111111111",
"0111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"0111111100111111111111111111110101010010011000001111111111111111111110010001010001111111111111111111111",
"0111111100111111111111111111110011010100000000110111111111111111111111111111111110010100000000001000000",
"0111111100111111111111111111111111111111000101000111111111111111111111111111111111111111111111111111111",
"0010011100000001111110001100011111111111111111111111111111111111111111111111111111000000001111010111101",
"0111111100111111111111111111111111111110010011001100011000011111111111111111111111111111111111111111111",
"0010011100000001111111101100010111010001111111111111111111111111111111111111111111111111111111111111111",
"0010101100000111111111111111111111111110001010110111111111111111111111111111111111111111111111111111111",
"0111111100111111111111111111111111111110000100011100010010011111111111111111111111111111111111111111111",
"0111111100111111111111111111111111111111111111111111111111111111111111111111111111000000000111010111101",
"0010101011100001111111101100011111111110010100101111111111111111111110010001110000100000000000000111011",
"0010001011000111111111111111110111010011111111111111111111111111111111111111111111000000001110000100001",
"0111111100111001111111101000011111111111111111111111111111110001001000010001010001111111111111111111111",
"0010001011100000000100001101111111111111000110000111111111100011000001111111111110100000001000010111101",
"0010011100000111111111111111110110010001111111111100001010111111111111111111111111000000000000000111011",
"0001111001100100000100010100000111010011111111111111111111111111111111111111111111111111111111111111111",
"0111111100111001111111101000011111111110000100011111111111111111111110010001010001111111111111111111111",
"0111111100111000001000001101111111111111000110000111111111111111111111111111111111111111111111111111111",
"0010011011000000001100001101111111111111111111111100000010111111111110010001110000000000001000010111101",
"0111111100111111111111111111111111111111000010101100011000011111111111111111111111111111111111111111111",
"0001111001100100000100010100000111010011111111111111111111111111111111111111111111111111111111111111111",
"0001001011100111111111111111111111111111111111111100010001111111111111111111111111111111111111111111111",
"0111111100111111111111111111111111111111111111111111111111110001001001111111111111111111111111111111111",
"0111111100111111111111111111111111111111111111111111111111111111111111111111111111000000010001010111101",
"0111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"0111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"0111111100111111111111111111111111111111111111111111111111111111111111111111111110000000010100110111101",
"0010001011100111111111111111111111111110001100100111111111111111111111111111111111111111111111111111111",
"0111111100111111111111111111110110010011111111111111111111111111111111111111111111111111111111111111111",
"0001010001001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"0000010001010100000100010100001111111111111111111111111111101111000001111111111111111111111111111111111",
"0111111100111001111111101100010110010000000100011111111111110001100001111111111111111111111111111111111",
"0010101011000000011101110000111111111111111111111100010110011111111111111111111110000000111111110100001",
"0111111100111001111111101100011111111111000101100111111111110001001000010001110001111111111111111111111",
"0111111100111000000100010000001111111111000010111100011000011111111111111111111110100000010001110111101",
"0111111100111100000100110100000110010101111111111100010000011111111111111111111111111111111111111111111",
"0010001011100111111111111111110110010011111111111111111111111111111110101111000001111111111111111111111",
"0010011011100111111111111111111111111110000100101111111111111111111111111111111111111111111111111111111",
"0111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"0111111100111111111111111111111111111111111111111111111111110001001001111111111111111111111111111111111",
"0111111100111111111111111111111111111111111111111111111111111111111111111111111110100000001000110111101",
"0111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"0001111001111100000011010100001111111111111111111111111111111111111111111111111111111111111111111111111",
"0010011001100100000011110100001111111111111111111111111111111111111111111111111111111111111111111111111",
"0001101011100111111111111111110110001111111111111111111111110001000111111111111111111111111111111111111",
"0111111100111111111111111111111111111111111111111111111111110001001001111111111111111111111111111111111",
"0111111100111111111111111111111111111111111111111111111111111111111111111111111110100000001001110111101",
"0111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"0010011001000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"0111111100111111111111111111111111111111111111111111111111111111111111111111111110000000000010010111101",
"0111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"0111111100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");

end snappy_tta_imem_image;
