library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use work.snappy_tta_imem_mau.all;

package snappy_tta_imem_image is

  type std_logic_imem_matrix is array (natural range <>) of std_logic_vector(IMEMMAUWIDTH-1 downto 0);

  constant imem_array : std_logic_imem_matrix := (
"0111111110111100000000000000001110111111111111111111111111111111111111111111111111110001111111111111111",
"1111111110111100000001001010100110111111111111111111111111111111111100000000000000000000000000000000011",
"0111111110111111000000000100111110111111111111111111111111111111111111111111111111110110000000001001100",
"0111111110111100000010001011100110111111100001101011111111111111111111111111111111100000000011100101100",
"0111111110111111111111111111111101000000010010000010001011001111111111111111111111111000000000001000100",
"0111111110111100000000001001100110111111111111111111111111111111111111111111111111111100000000001000100",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111100000000010010101100",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111100000000000000001110111111010011000011111111111111111111000000001101010001111111111111111",
"0111111110111111111111111111111101000000111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111100000000010110101101",
"0111111110111111111111111111111110111111111111111111111111110100100000000000010110010001111111111111111",
"0111111110111110000000011001100110111111111111111111111111111111111111111111111111111100000000001000100",
"0111111110111100000011110000101110111111111111111111111111111111111111111111111111100000000101010101101",
"0111111110111100000000010000100110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111100000000000000001110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111001100000111111111111111111110111111000111111111111100001000011100100101",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101011111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111100000110000110111110111111111111111111111111111111111111110000011000010001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111110000011000010001111111111111111",
"1111111110111100000100000110111101000110111111111111111111110000000000000000000001100000000111111000000",
"0111111110111111000000000100001110111111111111111110001010001111111111110000011000010001111111111111111",
"1111111110111100000010000110111110111111000010101111111111111100000000000000000000000000000000000111111",
"0111111110111111000000000100001110111111100001010110001010001111111111000011011000010001111111111111111",
"0111111110111100111111110100001110111111100011000010000101011111111111110000010100010001111111111111111",
"1111111110111111111111111111111110111111100011000010000101010000000000000111111110000000000000110000000",
"0111111110111111000000001101000101100000111111111111111111111111111111111111111111100000110000000100000",
"0111111110111111111111111111111101000110111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"1111111110111111111111111111111110111111111111111111111111110100011000000000001000000000000100010010011",
"0111111110111111111111111111111010110000111111111111111111111111111111000011011010000001011000110101001",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111100110000000110001011000110111111111111111111111111111111110000011000010001111111111111111",
"0111111110111100010000001101000101100000000010101111111111111111111111111111111111100000000101000101001",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111100000010000110001110111111111111111111111111111111111111000011011000010001111111111111111",
"0111111110111111111111111111111101100000000011100011111111111111111111111111111111100000001110010100000",
"0111111110111100000100000100001110111111111111111111111111111111111111000011010100010001111111111111111",
"0111111110111111111111111111111001000111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111100000000001001011110111111000011100011111111111111111111000011111010000000010000110101001",
"0111111110111111111111111111111110111111010001000111111111111111111111000011011000010001111111111111111",
"0111111110111111111111111111111101000110111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111100000100000110101101",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111110000010100010001111111111111111",
"0111111110111100111111110100001110111111111111111111111111111111111111110000011000010001111111111111111",
"1111111110111100000010000110111110111111000010101111111111111100000000000000000000000000000000000111111",
"0111111110111111000000000100001001000111111111111110001010001111111111111111111111110001111111111111111",
"0000111110010011111111111111111110111111000010101111111111111111111111110000011000011000000000000110101",
"1111111110111100000100000110111001000111111111111111111111110000000000000000000001100000000111111000000",
"0111111110111111000000000100001011001000111111111110001010001111111111110000011000010001111111111111111",
"1111111110111100000110000110111110111111111111111111111111110000000000000011111110000000000000000000000",
"0111111110111111000000000100001110111111100011000010001010001111111111000011101010110001111111111111111",
"0111111110111111111111111111111110111111100011000010000101011111111111111111111111110001111111111111111",
"0111111110111111111111111111111101100000000011100011111111111111111111111111111111100000111101000100000",
"0111111110111111111111111111111101000111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111000100000100110001111111111111111",
"0111111110111111111111111111111001100000000011100011111111111111111111111111111111100000011111110100111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111100000010110100101101",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0000001000100111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111110000010101100000110111111111111111111111111111111111111111111111111111100000000001001001",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111011001000010001100111111111111111111111110000011000010001111111111111111",
"0111111110111100000011110110001110111111111111111110001100001111111111111111111111110001111111111111111",
"0111111110111100000011111101000101100000111111111111111111111111111111111111111111100000011010000101001",
"0111111110111111111111111111111101001010000110000011111111111111111111000100110110010001111111111111111",
"0111111110111111111111111111111100001001111111111111111111111111111111111111111111110001111111111111111",
"0000101000101011111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111100111111110110001110111111111111111111111111111111111111110000011000010001111111111111111",
"0111111110111100111111111101000101100000000110000011111111111111111111000100110110000000011000100100000",
"0111111110111111111111111111111100001001111111111110001000001111111111000101010110010001111111111111111",
"0111111110111111111111111111111100001010111111111111111111111111111111111111111111110001111111111111111",
"0101010110011010100010101001000110111111111111111111111111111111111111000100110000010001111111111111111",
"0000111110110011111111111111111100100000000010101111111111111111111111111111111111100000001111110100010",
"0111111110111111111111111111111100001001111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111011001010111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0001010110010000111111110100001110111111111111111111111111111111111111110000011000010001111111111111111",
"1111111110111100000010000110111110111111111111111111111111111100000000000000000000000000000000000111111",
"0111111110111111000000000100001001001010001010000010001010001111111111000100110110010001111111111111111",
"0111111110111100000011110110001100001001111111111111111111111111111111000100011000010001111111111111111",
"0111111110111100000011111101000101100000111111111111111111111111111111111111111111100000010110010101001",
"0111111110111111111111111111111101001000100000010111111111111111111111000101010100010001111111111111111",
"0111111110111111111111111111111001001010010010000011111111111111111111000100010110010001111111111111111",
"0000101000100011111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111100111111110110001110111111111111111111111111111111111111110000011000010001111111111111111",
"0111111110111100111111111101000101100000000110000011111111111111111111000100110110000000011101100100000",
"0111111110111111111111111111111100001001111111111110001000001111111111000100010110010001111111111111111",
"0111111110111111111111111111111100001000111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111100000010110010101101",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111010010000011111111111111111111000100010110010001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111100000010000110101101",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0000111110000011111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0000111110000011111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111110000010100010001111111111111111",
"0111111110111100111111110100001110111111111111111111111111111111111111110000011000010001111111111111111",
"1111111110111100000010000110111110111111000010101111111111111100000000000000000000000000000000000111111",
"0111111110111111000000000100001001000111111111111110001010001111111111111111111111110001111111111111111",
"0000111110010011111111111111111110111111000010101111111111111111111111110000011000011000000000000110101",
"1111111110111100000100000110111001000111111111111111111111110000000000000000000001100000000111111000000",
"0111111110111111000000000100001011001000111111111110001010001111111111110000011000010001111111111111111",
"1111111110111100000110000110111110111111111111111111111111110000000000000011111110000000000000000000000",
"0111111110111111000000000100001110111111100011000010001010001111111111000011101010110001111111111111111",
"0111111110111111111111111111111110111111100011000010000101011111111111111111111111110001111111111111111",
"0111111110111111111111111111111101100000000011100011111111111111111111111111111111100000111101000100000",
"0111111110111111111111111111111101000111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111000100000100110001111111111111111",
"0111111110111111111111111111111001100000000011100011111111111111111111111111111111100000100000100100111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111100000100110100101101",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0000001000100111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111110000010101100000110111111111111111111111111111111111111111111111111111100000000001001001",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111011001000010001100111111111111111111111110000011000010001111111111111111",
"0111111110111100000011110110001110111111111111111110001100001111111111111111111111110001111111111111111",
"0111111110111100000011111101000101100000111111111111111111111111111111111111111111100000101010000101001",
"0111111110111111111111111111111101001010000110000011111111111111111111000100110110010001111111111111111",
"0111111110111111111111111111111100001001111111111111111111111111111111111111111111110001111111111111111",
"0000101000101011111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111100111111110110001110111111111111111111111111111111111111110000011000010001111111111111111",
"0111111110111100111111111101000101100000000110000011111111111111111111000100110110000000101000100100000",
"0111111110111111111111111111111100001001111111111110001000001111111111000101010110010001111111111111111",
"0111111110111111111111111111111100001010111111111111111111111111111111111111111111110001111111111111111",
"0101010110011011111111111111111110111111111111111111111111111111111111000100110000010001111111111111111",
"0111111110111111111111111111111100100000111111111111111111111111111111000011111100000000100000110100010",
"0111111110111111111111111111111100001001111111111111111111111111111111111111111111110001111111111111111",
"0001010110000011111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111110000010100010001111111111111111",
"0111111110111100111111110100001110111111111111111111111111111111111111110000011000010001111111111111111",
"1111111110111100000010000110111110111111111111111111111111111100000000000000000000000000000000000111111",
"0111111110111111000000000100001001001010001010000010001010001111111111000100110110010001111111111111111",
"0111111110111100000011110110001100001001111111111111111111111111111111000100011000010001111111111111111",
"0111111110111100000011111101000101100000111111111111111111111111111111111111111111100000100110010101001",
"0111111110111111111111111111111101001000100000010111111111111111111111000101010100010001111111111111111",
"0111111110111111111111111111111001001010010010000011111111111111111111000100010110010001111111111111111",
"0000101000100011111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111100111111110110001110111111111111111111111111111111111111110000011000010001111111111111111",
"0111111110111100111111111101000101100000000110000011111111111111111111000100110110000000101101110100000",
"0111111110111111111111111111111100001001111111111110001000001111111111000100010110010001111111111111111",
"0111111110111111111111111111111100001000111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111100000100110010101101",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111010010000011111111111111111111000100010110010001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111100000110000110111110111111111111111111111111111111111111110000011000010001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111110000011000010001111111111111111",
"1111111110111100000100000110111101000110111111111111111111110000000000000000000001100000000111111000000",
"0111111110111111000000000100001110111111111111111110001010001111111111110000011000010001111111111111111",
"1111111110111100000010000110111110111111000010101111111111111100000000000000000000000000000000000111111",
"0111111110111111000000000100001110111111100001010110001010001111111111000011011000010001111111111111111",
"0111111110111100111111110100001110111111100011000010000101011111111111110000010100010001111111111111111",
"1111111110111111111111111111111110111111100011000010000101010101010000000011100110100000000001110011000",
"0111111110111111000000001101000101100000111111111111111111111111111111111111111111100001011000110101001",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111110000011000010001111111111111111",
"0111111110111100111111110100001110111111111111111111111111111111111111110000010100010001111111111111111",
"1111111110111100000010000110111110111111111111111111111111111100000000000000000000000000000000000111111",
"0111111110111111000000000100001110111111100011000010001010001111111111111111111111110001111111111111111",
"1111111110111111111111111111111110111111100001010111111111110001011001000000000000000000000000000011100",
"0111111110111111000000001101000101100000111111111111111111111111111111111111111111100001011000110101001",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111011000111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111110000010100010001111111111111111",
"0111111110111100111111110100001110111111000010101111111111111111111111110000011000010001111111111111111",
"1111111110111100000010000110111110111111111111111111111111111100000000000000000000000000000000000111111",
"0111111110111111000000000100001001000110111111111110001010001111111111110000011000010001111111111111111",
"1111111110111100000100000110111110111111111111111111111111110000000000000000000001100000000111111000000",
"0111111110111111000000000100001110111111100001010110001010001111111111000011011000010001111111111111111",
"0111111110111111111111111111111110111111100011000010000101011111111111111111111111110001111111111111111",
"0111111110111111111111111111111101100000000011100011111111111111111111111111111111100000000101000100000",
"0111111110111111111111111111111101000110111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111100111111110110001110111111111111111111111111111111111111000011111000010001111111111111111",
"0111111110111100111111011101000101100000111111111111111111111111111111111111111111100000111111010100011",
"0111111110111111111111111111111101001000111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000011100011111111111111111111000100011010000001000101100100000",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000111100011111111111111111111000100011010000000000100010101001",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111000011100100110001111111111111111",
"0111111110111111111111111111111110111111000010101011111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111100000000101010101101",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0000110110000011111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000011100011111111111111111111000011011010000000000101000100000",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111100000000101010101101",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101011111111111111111111111111111111110001111111111111111",
"0111111110111100111111101101000110111111111111111111111111111111111111000100011010000001000011100100000",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111100111111111101000110111111111111111111111111111111111111000100011010000000000100010101001",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111000011100100110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111100000000101010101101",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101011111111111111111111111111111111110001111111111111111",
"0000001000011111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000110000011111111111111111111000011110110010001111111111111111",
"0111111110111111111111111111111100100000111111111111111111111111111111000011011100000001000100000101000",
"0111111110111111111111111111111100000111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000110000011111111111111111111000011110110010001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111100000000101000101101",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0000001000011111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0000001000011011111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111100111111110100001110111111111111111111111111111111111111000011110100010001111111111111111",
"0111111110111100011111110110001011001000100010110011111111111111111111110000011000010001111111111111111",
"0111111110111111111111111111111110111111100001011110001100001111111111111111111111110001111111111111111",
"0111111110111100100000000110001101001001111111111111111111111111111111000100011000010001111111111111111",
"0111111110111100000001111000000101100000000011100011111111111111111111111111111111100001000110110101001",
"0000110110011011111111111111111100000111111111111111111111111111111111010100110000010001111111111111111",
"0111111110111111111111111111111100000110111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000011100011111111111111111111000011011010000000000101000100000",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111100001001100100101101",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0000001000011111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111010101011110001100001111111111111111111111110001111111111111111",
"0101000011010111111111111111111110111111011101000110001010001111111111000100111000010001111111111111111",
"0111111110111111111111111111111001001010010010000010001011001111111111111111111111110001111111111111111",
"0111111110111111111111111111111100001000111111111111111111111111111111111111111111110001111111111111111",
"0001000110000110100010101100000110111111111111111111111111111111111111111111111111110001111111111111111",
"0100111110011011111111111111111110111111111111111111111111111111111111000100010000010001111111111111111",
"0111111110111111111111111111111100100000111111111111111111111111111111000011011100000000000101000100010",
"0111111110111111111111111111111100000111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111110000011000010001111111111111111",
"0111111110111100111111000100001011001000111111111111111111111111111111110000010100010001111111111111111",
"0111111110111111111111111111111001001001001101000111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111101100000000011100011111111111111111111111111111111100001010011100100000",
"0111111110111111111111111111111101001011001001100111111111111111111111000100111000010001111111111111111",
"0111111110111100111111110110001101001001111111111111111111111111111111000100011000010001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000111100011111111111111111111000101111010000001001010010100000",
"0111111110111100111111110110001110111111111111111111111111111111111111110000011000010001111111111111111",
"0111111110111100001110000110001101001000111111111111111111111111111111000100111000010001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111110000011000010001111111111111111",
"1111111110111100000010000110111110111111111111111111111111111100000000000000000000000000000000000111111",
"0111111110111111000000000110001110111111111111111110001100001111111111111111111111110001111111111111111",
"0101000110100011111111111111111110111111001011100010000101011111111111000101111010000001001011010100000",
"0111111110111111111111111111111101001010000110000011111111111111111111000100110110010001111111111111111",
"0111111110111111111111111111111100001000111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111110000011000010001111111111111111",
"1111111110111100000100000110111110111111000010101111111111110000000000000000000001100000000111111000000",
"0111111110111111000000000100001110111111111111111110001010001111111111111111111111110001111111111111111",
"0001010110010000000110000110111110111111100000010111111111111111111111110000011000000001001011010101101",
"0111111110111111111111111111111110111111100001010110001100001111111111111111111111110001111111111111111",
"0111111110111111111111111111111101001010111111111111111111111111111111111111111111110001111111111111111",
"0111111110111100111100001101000101100000111111111111111111111111111111111111111111100001010101000100010",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111100001001011100101101",
"0111111110111111111111111111111110111111000110000011111111111111111111000100110110010001111111111111111",
"0111111110111111111111111111111100001000111111111111111111111111111111111111111111111100000000001001000",
"0000100000100011111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0000001000101011111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111100111111110110001110111111111111111111111111111111111111110000011000010001111111111111111",
"0111111110111100111111110100001110111111111111111111111111111111111111000101010100010001111111111111111",
"0111111110111100000010001000000101001011100010110011111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111100001010111111111111111111110111100000000100110110010001111111111111111",
"0111111110111100111111110110001100001001111111111111111111111000110000111111111111110001111111111111111",
"0111111110111100001110111101000101100000100001011111111111111111111111000101111000000001010101100100100",
"0001000110011011111111111111111110111111111111111110001000001111111111111111111111110001111111111111111",
"0111111110111111111111111111111100001000111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111100001001011110101101",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0001000110000010100001111011000110111111111111111111111111111111111111000100010000010001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110110000000000101101",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111100000000010000001110111111111111111111111111111111111111111111111111110001111111111111111");

end snappy_tta_imem_image;
