library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use work.snappy_tta_imem_mau.all;

package snappy_tta_imem_image is

  type std_logic_imem_matrix is array (natural range <>) of std_logic_vector(IMEMMAUWIDTH-1 downto 0);

  constant imem_array : std_logic_imem_matrix := (
"0111111110111100000000000000001110111111111111111111111111111111111111111111111111110001111111111111111",
"1111111110111100000001001010100110111111111111111111111111111111111100000000000000000000000000000000011",
"0111111110111111000000000100111110111111111111111111111111111111111111111111111111110110000000001001100",
"0111111110111100000010001011100110111111100001101011111111111111111111111111111111100000000001100101100",
"0111111110111111111111111111111101000000010010000010001011001111111111111111111111111000000000001000100",
"0111111110111100000000001001100110111111111111111111111111111111111111111111111111111100000000001000100",
"0111111110111100001110110000110110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111100000000010000101110111111111111111111111111111111111111111111111111100000000010110101101",
"0111111110111100111100000000100110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111100000000000000001110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101011111111111111111111111111111111110001111111111111111",
"0000001000011111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0000001000100011111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111100111111110100001110111111111111111111111111111111111111000100010100010001111111111111111",
"0111111110111100011111110110001011001001100010110011111111111111111111110000011000010001111111111111111",
"0111111110111111111111111111111110111111100001011110001100001111111111111111111111110001111111111111111",
"0111111110111100100000000110001101001010111111111111111111111111111111000100111000010001111111111111111",
"0111111110111111111111111111111101100000011110000011111111111111111111000000111100000000000011010101001",
"0000111110011011111111111111111100001000111111111111111111111111111111010101010000010001111111111111111",
"0111111110111111111111111111111100000111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000011100011111111111111111111000011111010000000000010100100000",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111100000001001000101101",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0000001000100011111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111010101011110001100001111111111111111111111110001111111111111111",
"0101001011010111111111111111111110111111011101000110001010001111111111000101011000010001111111111111111",
"0111111110111111111111111111111001001011010010000010001011001111111111111111111111110001111111111111111",
"0111111110111111111111111111111100001001111111111111111111111111111111111111111111110001111111111111111",
"0001001110000110100010111100000110111111111111111111111111111111111111111111111111110001111111111111111",
"0101000110011011111111111111111110111111111111111111111111111111111111000100110000010001111111111111111",
"0111111110111111111111111111111100100000111111111111111111111111111111000011111100000000000010100100010",
"0111111110111111111111111111111100001000111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111100111111000100001011001001001101000111111111111111111111110000011000011010000000001010100",
"0111111110111111111111111111111101100000100011000011111111111111111111000000111100000000001111100100000",
"0111111110111111111111111111111101001100001001100111111111111111111111111111111111110001111111111111111",
"0111111110111100111111110110001101001010111111111111111111111111111111000100111000010001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0100101110110011111111111111111110111111111111111111111111111111111111000110011010000000000110110100000",
"0111111110111100111111110110001110111111111111111111111111111111111111110000011000010001111111111111111",
"0111111110111100001110000110001101001001111111111111111111111111111111000101011000010001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111110000011000010001111111111111111",
"1111111110111100000010000110111110111111111111111111111111111100000000000000000000000000000000000111111",
"0111111110111111000000000110001110111111111111111110001100001111111111111111111111110001111111111111111",
"0101001110100011111111111111111110111111001011100010000101011111111111000110011010000000000111110100000",
"0111111110111111111111111111111101001011000110000011111111111111111111000101010110010001111111111111111",
"0111111110111111111111111111111100001001111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111110000011000010001111111111111111",
"1111111110111100000100000110111110111111000010101111111111110000000000000000000001100000000111111000000",
"0111111110111111000000000100001110111111111111111110001010001111111111111111111111110001111111111111111",
"0001011110010000000110000110111110111111100000010111111111111111111111110000011000000000000111110101101",
"0111111110111111111111111111111110111111100001010110001100001111111111111111111111110001111111111111111",
"0111111110111111111111111111111101001011111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111101100000111111111111111111111111111111000010011100000000010001000100010",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111100000001000000101101",
"0111111110111111111111111111111110111111000110000011111111111111111111000101010110010001111111111111111",
"0111111110111111111111111111111100001001111111111111111111111111111111111111111111111100000000001001000",
"0000101000100111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0000001000101111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111100111111110110001110111111111111111111111111111111111111000101111000010001111111111111111",
"0111111110111100111111110100001110111111111111111111111111111111111111110000010100010001111111111111111",
"0111111110111111111111111111111101001011100011000010000101111111111111111111111111110001111111111111111",
"0111111110111111111111111111111101001100111111111111111111110111100000000101010110010001111111111111111",
"0111111110111100111111110110001100001010111111111111111111111000110000111111111111110001111111111111111",
"0101011110011000000010001000000101100000111111111111111111111111111111000011011100000000010001100100100",
"0001001110011011111111111111111100001011111111111111111111111111111111010110010000010001111111111111111",
"0111111110111111111111111111111100001001111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111100000001000010101101",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0001001110000010100010001011000110111111111111111111111111111111111111000100110000010001111111111111111");

end snappy_tta_imem_image;
