library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use work.snappy_tta_imem_mau.all;

package snappy_tta_imem_image is

  type std_logic_imem_matrix is array (natural range <>) of std_logic_vector(IMEMMAUWIDTH-1 downto 0);

  constant imem_array : std_logic_imem_matrix := (
"0111111110111100000000000000001110111111111111111111111111111111111111111111111111110001111111111111111",
"1111111110111100000001001010100110111111111111111111111111111111111100000000000000000000000000000000011",
"0111111110111111000000000100111110111111111111111111111111111111111111111111111111110110000000001001100",
"0111111110111100000010001011100110111111100001101011111111111111111111111111111111100000000011010101100",
"0111111110111111111111111111111101000000010010000010001011001111111111111111111111111000000000001000100",
"0111111110111100000000001001100110111111111111111111111111111111111111111111111111111100000000001000100",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111100000000010010101100",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111100000001000000001110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111100000000010100101101",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0000001101010000000000001001100110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111100000011110001110110111111111111111111111111111111111111111111111111110001111111111111111",
"1111111110111100010000000001101110111111111111111111111111110100011000000000001000000000000100010010011",
"0111111110111111111111111111111010001100111111111111111111111111111111111111111111110001111111111111111",
"0111111110111100111111110001011110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111101111111110001010110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111100001110110001001110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111100000000010001000110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111100111100000000111110111111111111111111111111111111111111111111111111110001111111111111111",
"1111111110111100000000000000110110111111111111111111111111110001011001000000000000000000000000000011100",
"0111111110111100111111010000101110111111111111111111111111111111111111111111111111100000000110100101101",
"1111111110111111111111111111111010000100111111111111111111110101010000000011100110100000000001110011000",
"0111111110111111111111111111111010000001111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101011111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111100000110000110111110111111111111111111111111111111111111110000011000010001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111110000011000010001111111111111111",
"1111111110111100000100000110111101001111111111111111111111110000000000000000000001100000000111111000000",
"0111111110111111000000000100001110111111111111111110001010001111111111110000011000010001111111111111111",
"1111111110111100000010000110111110111111000010101111111111111100000000000000000000000000000000000111111",
"0111111110111111000000000100001110111111100001010110001010001111111111000111111000010001111111111111111",
"0111111110111100111111110100001110111111100011000010000101011111111111110000010100010001111111111111111",
"1111111110111111111111111111111110111111100011000010000101010000000000000111111110000000000000110000000",
"0111111110111111000000001101000101100000111111111111111111111111111111111111111111100000110001000100000",
"0111111110111111111111111111111101001111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0101100110110011111111111111111110111111111111111111111111111111111111000111111010000001011011000101001",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111100110000000110001011010000111111111111111111111111111111110000011000010001111111111111111",
"0111111110111111111111111111111101100000000010101111111111111111111111000110111100000000000110010101001",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111100000010000110001110111111111111111111111111111111111111001000011000010001111111111111111",
"0111111110111111111111111111111101100000000011100011111111111111111111111111111111100000001111010100000",
"0111111110111100000100000100001110111111111111111111111111111111111111001000010100010001111111111111111",
"0111111110111111111111111111111001001111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111100000000001001011110111111000011100011111111111111111111000111111010000000010001110101001",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111100000100001100101101",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111110000010100010001111111111111111",
"0111111110111100111111110100001110111111111111111111111111111111111111110000011000010001111111111111111",
"1111111110111100000010000110111110111111000010101111111111111100000000000000000000000000000000000111111",
"0111111110111111000000000100001001001111111111111110001010001111111111111111111111110001111111111111111",
"0001111110010011111111111111111110111111000010101111111111111111111111110000011000011000000000000110101",
"1111111110111100000100000110111001001111111111111111111111110000000000000000000001100000000111111000000",
"0111111110111111000000000100001011010000111111111110001010001111111111110000011000010001111111111111111",
"1111111110111100000110000110111110111111111111111111111111110000000000000011111110000000000000000000000",
"0111111110111111000000000100001110111111100011000010001010001111111111000111101010110001111111111111111",
"0111111110111111111111111111111110111111100011000010000101011111111111111111111111110001111111111111111",
"0111111110111111111111111111111101100000000011100011111111111111111111111111111111100000000110010100000",
"0111111110111111111111111111111101001111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111001000000100110001111111111111111",
"0111111110111111111111111111111001100000111111111111111111111111111111000011011100000000100000100100111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111100000010111100101101",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0000110001000011111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111110000100101100000110111111111111111111111111111111111111111111111111111100000000001001001",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111100111100000110001011010001111111111111111111111111111111110000011000010001111111111111111",
"0111111110111111111111111111111101100000111111111111111111111111111111000011111100000000011010100101001",
"0111111110111111111111111111111110111111000110000011111111111111111111001000010110010001111111111111111",
"0111111110111111111111111111111100010000111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111100111111110110001110111111111111111111111111111111111111110000011000010001111111111111111",
"0111111110111100111111111101000101100000111111111111111111111111111111111111111111100000011001000100000",
"0111111110111111111111111111111110111111000110000011111111111111111111001000010110010001111111111111111",
"0111111110111111111111111111111100010000111111111111111111111111111111111111111111110001111111111111111",
"0101111110011010100011111001000110111111111111111111111111111111111111001000010000010001111111111111111",
"0111111110111111111111111111111100100000000010101111111111111111111111001000011100000000010000110100010",
"0111111110111111111111111111111100010011111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111011010010111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0010010110010000111111110100001110111111111111111111111111111111111111110000011000010001111111111111111",
"1111111110111100000010000110111110111111111111111111111111111100000000000000000000000000000000000111111",
"0111111110111111000000000100001001010000111111111110001010001111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111100000010111111111111111111111001000010100010001111111111111111",
"0111111110111100000011110110001001010010111111111111111111111111111111001000111000010001111111111111111",
"0111111110111111111111111111111101100000111111111111111111111111111111000111011100000000010111010101001",
"0111111110111111111111111111111101010001001010000011111111111111111111001001110110010001111111111111111",
"0111111110111111111111111111111100010000010010000011111111111111111111001000110110010001111111111111111",
"0001110001000111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111100111111110110001110111111111111111111111111111111111111110000011000010001111111111111111",
"0111111110111100111111111101000101100000000110000011111111111111111111001000010110000000011110010100000",
"0111111110111111111111111111111100010000111111111110001000001111111111001000110110010001111111111111111",
"0111111110111111111111111111111100010001111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111100000010111010101101",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111010010000011111111111111111111001000110110010001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111100000010001110101101",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0001111110000011111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0001111110000011111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111110000010100010001111111111111111",
"0111111110111100111111110100001110111111111111111111111111111111111111110000011000010001111111111111111",
"1111111110111100000010000110111110111111000010101111111111111100000000000000000000000000000000000111111",
"0111111110111111000000000100001001001111111111111110001010001111111111111111111111110001111111111111111",
"0001111110010011111111111111111110111111000010101111111111111111111111110000011000011000000000000110101",
"1111111110111100000100000110111001001111111111111111111111110000000000000000000001100000000111111000000",
"0111111110111111000000000100001011010000111111111110001010001111111111110000011000010001111111111111111",
"1111111110111100000110000110111110111111111111111111111111110000000000000011111110000000000000000000000",
"0111111110111111000000000100001110111111100011000010001010001111111111000111101010110001111111111111111",
"0111111110111111111111111111111110111111100011000010000101011111111111111111111111110001111111111111111",
"0111111110111111111111111111111101100000000011100011111111111111111111111111111111100000000110010100000",
"0111111110111111111111111111111101001111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111001000000100110001111111111111111",
"0111111110111111111111111111111001100000111111111111111111111111111111000011011100000000100001010100111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111100000100111010101101",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0000110001000011111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111110000100101100000110111111111111111111111111111111111111111111111111111100000000001001001",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111100111100000110001011010001111111111111111111111111111111110000011000010001111111111111111",
"0111111110111111111111111111111101100000111111111111111111111111111111000011111100000000101010010101001",
"0111111110111111111111111111111110111111000110000011111111111111111111001000010110010001111111111111111",
"0111111110111111111111111111111100010000111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111100111111110110001110111111111111111111111111111111111111110000011000010001111111111111111",
"0111111110111100111111111101000101100000111111111111111111111111111111111111111111100000101000110100000",
"0111111110111111111111111111111110111111000110000011111111111111111111001000010110010001111111111111111",
"0111111110111111111111111111111100010000111111111111111111111111111111111111111111110001111111111111111",
"0101111110011011111111111111111110111111111111111111111111111111111111001000010000010001111111111111111",
"0111111110111111111111111111111100010011111111111111111111111000100011001000010110010001111111111111111",
"0111111110111111111111111111111110111111000100101011111111111000101000111111111111110001111111111111111",
"0111111110111111111111111111111001100000111111111111111111111111111111111111111111100000100001100101010",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0001111110000011111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111110000010100010001111111111111111",
"0111111110111100111111110100001110111111111111111111111111111111111111110000011000010001111111111111111",
"1111111110111100000010000110111110111111111111111111111111111100000000000000000000000000000000000111111",
"0111111110111111000000000100001001010000111111111110001010001111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111100000010111111111111111111111001000010100010001111111111111111",
"0111111110111100000011110110001001010010111111111111111111111111111111001000111000010001111111111111111",
"0111111110111111111111111111111101100000111111111111111111111111111111000111011100000000100111000101001",
"0111111110111111111111111111111101010001001010000011111111111111111111001001110110010001111111111111111",
"0111111110111111111111111111111100010000010010000011111111111111111111001000110110010001111111111111111",
"0001110001000111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111100111111110110001110111111111111111111111111111111111111110000011000010001111111111111111",
"0111111110111100111111111101000101100000000110000011111111111111111111001000010110000000101110110100000",
"0111111110111111111111111111111100010000111111111110001000001111111111001000110110010001111111111111111",
"0111111110111111111111111111111100010001111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111100000100111000101101",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111010010000011111111111111111111001000110110010001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111100000110000110111110111111111111111111111111111111111111110000011000010001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111110000011000010001111111111111111",
"1111111110111100000100000110111101001111111111111111111111110000000000000000000001100000000111111000000",
"0111111110111111000000000100001110111111111111111110001010001111111111110000011000010001111111111111111",
"1111111110111100000010000110111110111111000010101111111111111100000000000000000000000000000000000111111",
"0111111110111111000000000100001110111111100001010110001010001111111111000111111000010001111111111111111",
"0111111110111100111111110100001110111111100011000010000101011111111111110000010100010001111111111111111",
"0111111110111111111111111111111110111111100011000010000101011111111111111111111111110001111111111111111",
"0111111110111111111111111111111101100000111111111111111111111111111111000000111100000001011011000101001",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111110000011000010001111111111111111",
"0111111110111100111111110100001110111111111111111111111111111111111111110000010100010001111111111111111",
"1111111110111100000010000110111110111111111111111111111111111100000000000000000000000000000000000111111",
"0111111110111111000000000100001110111111100011000010001010001111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111100001010111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111101100000111111111111111111111111111111000010011100000001011011000101001",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111011001111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111110000010100010001111111111111111",
"0111111110111100111111110100001110111111000010101111111111111111111111110000011000010001111111111111111",
"1111111110111100000010000110111110111111111111111111111111111100000000000000000000000000000000000111111",
"0111111110111111000000000100001001010000111111111110001010001111111111110000011000010001111111111111111",
"1111111110111100000100000110111110111111111111111111111111110000000000000000000001100000000111111000000",
"0111111110111111000000000100001110111111100001010110001010001111111111001000011000010001111111111111111",
"0111111110111111111111111111111110111111100011000010000101011111111111111111111111110001111111111111111",
"0111111110111111111111111111111101100000000011100011111111111111111111111111111111100001000001000101001",
"0111111110111111111111111111111101010000111111111111111111111111111111111111111111110001111111111111111",
"0111111110111100111111110110001110111111111111111111111111111111111111000111111000010001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111100000000110010101101",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000011100011111111111111111111001000111010000001000110000100000",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000111100011111111111111111111001000111010000001011000100101001",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111000111100100110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0010000110000011111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111011001111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111110000010100010001111111111111111",
"0111111110111100111111110100001110111111000010101111111111111111111111110000011000010001111111111111111",
"1111111110111100000010000110111110111111111111111111111111111100000000000000000000000000000000000111111",
"0111111110111111000000000100001001010000111111111110001010001111111111110000011000010001111111111111111",
"1111111110111100000100000110111110111111111111111111111111110000000000000000000001100000000111111000000",
"0111111110111111000000000100001110111111100001010110001010001111111111001000011000010001111111111111111",
"0111111110111111111111111111111110111111100011000010000101011111111111111111111111110001111111111111111",
"0111111110111111111111111111111101100000111111111111111111111111111111000011011100000000000110010100000",
"0111111110111111111111111111111101010000111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111100111111110110001110111111111111111111111111111111111111000111111000010001111111111111111",
"0111111110111111111111111111111101100000111111111111111111111111111111000010111100000000111010110100101",
"0111111110111111111111111111111101010001111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111100111111101101000110111111111111111111111111111111111111001000111010000001011001100100000",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111110111100000001000010110010001111111111111111",
"0101011110110011111111111111111110111111111111111111111111111111111111001000111010000001011000100101001",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111000111100100110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111100000111101100101101",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0000110001000011111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0000110000111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111100111111110100001110111111111111111111111111111111111111001000010100010001111111111111111",
"0111111110111100011111110110001011010001100010110011111111111111111111110000011000010001111111111111111",
"0111111110111111111111111111111110111111100001011110001100001111111111111111111111110001111111111111111",
"0111111110111100100000000110001101010010111111111111111111111111111111001000111000010001111111111111111",
"0111111110111111111111111111111101100000011110000011111111111111111111000011011100000001000111010101001",
"0001111110011011111111111111111100010000111111111111111111111111111111011001010000010001111111111111111",
"0111111110111111111111111111111100001111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000011100011111111111111111111000111111010000000111101100100000",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111100001001101000101101",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0000110001000011111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111010101011110001100001111111111111111111111110001111111111111111",
"0110001011010111111111111111111110111111011101000110001010001111111111001001011000010001111111111111111",
"0111111110111111111111111111111001010011010010000010001011001111111111111111111111110001111111111111111",
"0111111110111111111111111111111100010001111111111111111111111111111111111111111111110001111111111111111",
"0010001110000110100100111100000110111111111111111111111111111111111111111111111111110001111111111111111",
"0110000110011011111111111111111110111111111111111111111111111111111111001000110000010001111111111111111",
"0111111110111111111111111111111100100000111111111111111111111111111111000111111100000000111101100100010",
"0111111110111111111111111111111100010000111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111100111111000100001011010001001101000111111111111111111111110000011000011010000000001010100",
"0111111110111111111111111111111101100000100011000011111111111111111111000011011100000001010011100100000",
"0111111110111111111111111111111101010100001001100111111111111111111111111111111111110001111111111111111",
"0111111110111100111111110110001101010010111111111111111111111111111111001000111000010001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0101000110110011111111111111111110111111111111111111111111111111111111001010011010000001001010110100000",
"0111111110111100111111110110001110111111111111111111111111111111111111110000011000010001111111111111111",
"0111111110111100001110000110001101010001111111111111111111111111111111001001011000010001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111110000011000010001111111111111111",
"1111111110111100000010000110111110111111111111111111111111111100000000000000000000000000000000000111111",
"0111111110111111000000000110001110111111111111111110001100001111111111111111111111110001111111111111111",
"0110001110100011111111111111111110111111001011100010000101011111111111001010011010000001001011110100000",
"0111111110111111111111111111111101010011000110000011111111111111111111001001010110010001111111111111111",
"0111111110111111111111111111111100010001111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111110000011000010001111111111111111",
"1111111110111100000100000110111110111111000010101111111111110000000000000000000001100000000111111000000",
"0111111110111111000000000100001110111111111111111110001010001111111111111111111111110001111111111111111",
"0010011110010000000110000110111110111111100000010111111111111111111111110000011000000001001011110101101",
"0111111110111111111111111111111110111111100001010110001100001111111111111111111111110001111111111111111",
"0111111110111111111111111111111101010011111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111101100000111111111111111111111111111111000011111100000001010101000100010",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111100001001100000101101",
"0111111110111111111111111111111110111111000110000011111111111111111111001001010110010001111111111111111",
"0111111110111111111111111111111100010001111111111111111111111111111111111111111111111100000000001001000",
"0001000001000111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0000110001001111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111000010101111111111111111111111111111111111110001111111111111111",
"0111111110111100111111110110001110111111111111111111111111111111111111001001111000010001111111111111111",
"0111111110111100111111110100001110111111111111111111111111111111111111110000010100010001111111111111111",
"0111111110111111111111111111111101010011100011000010000101111111111111111111111111110001111111111111111",
"0111111110111111111111111111111101010100111111111111111111110111100000001001010110010001111111111111111",
"0111111110111100111111110110001100010010111111111111111111111000110000111111111111110001111111111111111",
"0110011110011000000010001000000101100000111111111111111111111111111111000100111100000001010101100100100",
"0010001110011011111111111111111100010011111111111111111111111111111111011010010000010001111111111111111",
"0111111110111111111111111111111100010001111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111100001001100010101101",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0010001110000010100100001011000110111111111111111111111111111111111111001000110000010001111111111111111",
"0111111110111111111111111111111001100000111111111111111111111111111111000101011100000000000110010100110",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111110111100000001000010110010001111111111111111",
"0111111110111111111111111111111100100000111111111111111111111111111111000011011100000001011001100101001",
"0111111110111111111111111111111100010000000010101111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111110111100000001000010110010001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111100000111101100101101",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110110000000000101101",
"0111111110111111111111111111111110111111111111111111111111111111111111111111111111110001111111111111111",
"0111111110111100000000010000001110111111111111111111111111111111111111111111111111110001111111111111111");

end snappy_tta_imem_image;
