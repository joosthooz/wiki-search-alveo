package snappy_tta_params is
  constant fu_LSU_addrw_g : integer := 12;
end snappy_tta_params;
