package snappy_tta_imem_mau is
   -- created by generatebits
   constant IMEMMAUWIDTH : positive := 107;
end snappy_tta_imem_mau;
